library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity jalfunction is
	port (x: in std_logic);
end jalfunction;

architecture beh of jalfunction is
begin
end beh;
